********************************************************************************
* Revolution EDA CDL Netlist
* Library: designs
* Top Cell Name: lowPassFilter
* View Name: schematic
* Date: 2022-07-07 17:28:38.884588
********************************************************************************
.GLOBAL gnd!

XI2 INP net0 lowPassRC
XI3 net0 OUT lowPassRC
.END
